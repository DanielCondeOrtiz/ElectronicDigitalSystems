LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

--Declaraci�n de la entidad
ENTITY testa IS
END    testa;

ARCHITECTURE testa_arq OF testa IS
BEGIN


END testa_arq;












